----------------------------------------------------------------------------------
-- Module Name: SBox - SBox_architecture
-- Project Name: AES - Advanced Encryption Standard 
-- Description: Rijndael substitution box used in key expansion and cipher rounds.
----------------------------------------------------------------------------------

library IEEE;
use IEEE.STD_LOGIC_1164.ALL;

entity SBox is
port (
	INPUT  : in std_logic_vector(7 downto 0);   -- input byte
	OUTPUT : out std_logic_vector(7 downto 0)); -- output byte
end SBox;

architecture SBox_architecture of SBox is
begin
    process(INPUT)
    begin
        case INPUT is
            when "00000000" => OUTPUT <= "01100011";
            when "00000001" => OUTPUT <= "01111100";
            when "00000010" => OUTPUT <= "01110111";
            when "00000011" => OUTPUT <= "01111011";
            when "00000100" => OUTPUT <= "11110010";
            when "00000101" => OUTPUT <= "01101011";
            when "00000110" => OUTPUT <= "01101111";
            when "00000111" => OUTPUT <= "11000101";
            when "00001000" => OUTPUT <= "00110000";
            when "00001001" => OUTPUT <= "00000001";
            when "00001010" => OUTPUT <= "01100111";
            when "00001011" => OUTPUT <= "00101011";
            when "00001100" => OUTPUT <= "11111110";
            when "00001101" => OUTPUT <= "11010111";
            when "00001110" => OUTPUT <= "10101011";
            when "00001111" => OUTPUT <= "01110110";
            when "00010000" => OUTPUT <= "11001010";
            when "00010001" => OUTPUT <= "10000010";
            when "00010010" => OUTPUT <= "11001001";
            when "00010011" => OUTPUT <= "01111101";
            when "00010100" => OUTPUT <= "11111010";
            when "00010101" => OUTPUT <= "01011001";
            when "00010110" => OUTPUT <= "01000111";
            when "00010111" => OUTPUT <= "11110000";
            when "00011000" => OUTPUT <= "10101101";
            when "00011001" => OUTPUT <= "11010100";
            when "00011010" => OUTPUT <= "10100010";
            when "00011011" => OUTPUT <= "10101111";
            when "00011100" => OUTPUT <= "10011100";
            when "00011101" => OUTPUT <= "10100100";
            when "00011110" => OUTPUT <= "01110010";
            when "00011111" => OUTPUT <= "11000000";
            when "00100000" => OUTPUT <= "10110111";
            when "00100001" => OUTPUT <= "11111101";
            when "00100010" => OUTPUT <= "10010011";
            when "00100011" => OUTPUT <= "00100110";
            when "00100100" => OUTPUT <= "00110110";
            when "00100101" => OUTPUT <= "00111111";
            when "00100110" => OUTPUT <= "11110111";
            when "00100111" => OUTPUT <= "11001100";
            when "00101000" => OUTPUT <= "00110100";
            when "00101001" => OUTPUT <= "10100101";
            when "00101010" => OUTPUT <= "11100101";
            when "00101011" => OUTPUT <= "11110001";
            when "00101100" => OUTPUT <= "01110001";
            when "00101101" => OUTPUT <= "11011000";
            when "00101110" => OUTPUT <= "00110001";
            when "00101111" => OUTPUT <= "00010101";
            when "00110000" => OUTPUT <= "00000100";
            when "00110001" => OUTPUT <= "11000111";
            when "00110010" => OUTPUT <= "00100011";
            when "00110011" => OUTPUT <= "11000011";
            when "00110100" => OUTPUT <= "00011000";
            when "00110101" => OUTPUT <= "10010110";
            when "00110110" => OUTPUT <= "00000101";
            when "00110111" => OUTPUT <= "10011010";
            when "00111000" => OUTPUT <= "00000111";
            when "00111001" => OUTPUT <= "00010010";
            when "00111010" => OUTPUT <= "10000000";
            when "00111011" => OUTPUT <= "11100010";
            when "00111100" => OUTPUT <= "11101011";
            when "00111101" => OUTPUT <= "00100111";
            when "00111110" => OUTPUT <= "10110010";
            when "00111111" => OUTPUT <= "01110101";
            when "01000000" => OUTPUT <= "00001001";
            when "01000001" => OUTPUT <= "10000011";
            when "01000010" => OUTPUT <= "00101100";
            when "01000011" => OUTPUT <= "00011010";
            when "01000100" => OUTPUT <= "00011011";
            when "01000101" => OUTPUT <= "01101110";
            when "01000110" => OUTPUT <= "01011010";
            when "01000111" => OUTPUT <= "10100000";
            when "01001000" => OUTPUT <= "01010010";
            when "01001001" => OUTPUT <= "00111011";
            when "01001010" => OUTPUT <= "11010110";
            when "01001011" => OUTPUT <= "10110011";
            when "01001100" => OUTPUT <= "00101001";
            when "01001101" => OUTPUT <= "11100011";
            when "01001110" => OUTPUT <= "00101111";
            when "01001111" => OUTPUT <= "10000100";
            when "01010000" => OUTPUT <= "01010011";
            when "01010001" => OUTPUT <= "11010001";
            when "01010010" => OUTPUT <= "00000000";
            when "01010011" => OUTPUT <= "11101101";
            when "01010100" => OUTPUT <= "00100000";
            when "01010101" => OUTPUT <= "11111100";
            when "01010110" => OUTPUT <= "10110001";
            when "01010111" => OUTPUT <= "01011011";
            when "01011000" => OUTPUT <= "01101010";
            when "01011001" => OUTPUT <= "11001011";
            when "01011010" => OUTPUT <= "10111110";
            when "01011011" => OUTPUT <= "00111001";
            when "01011100" => OUTPUT <= "01001010";
            when "01011101" => OUTPUT <= "01001100";
            when "01011110" => OUTPUT <= "01011000";
            when "01011111" => OUTPUT <= "11001111";
            when "01100000" => OUTPUT <= "11010000";
            when "01100001" => OUTPUT <= "11101111";
            when "01100010" => OUTPUT <= "10101010";
            when "01100011" => OUTPUT <= "11111011";
            when "01100100" => OUTPUT <= "01000011";
            when "01100101" => OUTPUT <= "01001101";
            when "01100110" => OUTPUT <= "00110011";
            when "01100111" => OUTPUT <= "10000101";
            when "01101000" => OUTPUT <= "01000101";
            when "01101001" => OUTPUT <= "11111001";
            when "01101010" => OUTPUT <= "00000010";
            when "01101011" => OUTPUT <= "01111111";
            when "01101100" => OUTPUT <= "01010000";
            when "01101101" => OUTPUT <= "00111100";
            when "01101110" => OUTPUT <= "10011111";
            when "01101111" => OUTPUT <= "10101000";
            when "01110000" => OUTPUT <= "01010001";
            when "01110001" => OUTPUT <= "10100011";
            when "01110010" => OUTPUT <= "01000000";
            when "01110011" => OUTPUT <= "10001111";
            when "01110100" => OUTPUT <= "10010010";
            when "01110101" => OUTPUT <= "10011101";
            when "01110110" => OUTPUT <= "00111000";
            when "01110111" => OUTPUT <= "11110101";
            when "01111000" => OUTPUT <= "10111100";
            when "01111001" => OUTPUT <= "10110110";
            when "01111010" => OUTPUT <= "11011010";
            when "01111011" => OUTPUT <= "00100001";
            when "01111100" => OUTPUT <= "00010000";
            when "01111101" => OUTPUT <= "11111111";
            when "01111110" => OUTPUT <= "11110011";
            when "01111111" => OUTPUT <= "11010010";
            when "10000000" => OUTPUT <= "11001101";
            when "10000001" => OUTPUT <= "00001100";
            when "10000010" => OUTPUT <= "00010011";
            when "10000011" => OUTPUT <= "11101100";
            when "10000100" => OUTPUT <= "01011111";
            when "10000101" => OUTPUT <= "10010111";
            when "10000110" => OUTPUT <= "01000100";
            when "10000111" => OUTPUT <= "00010111";
            when "10001000" => OUTPUT <= "11000100";
            when "10001001" => OUTPUT <= "10100111";
            when "10001010" => OUTPUT <= "01111110";
            when "10001011" => OUTPUT <= "00111101";
            when "10001100" => OUTPUT <= "01100100";
            when "10001101" => OUTPUT <= "01011101";
            when "10001110" => OUTPUT <= "00011001";
            when "10001111" => OUTPUT <= "01110011";
            when "10010000" => OUTPUT <= "01100000";
            when "10010001" => OUTPUT <= "10000001";
            when "10010010" => OUTPUT <= "01001111";
            when "10010011" => OUTPUT <= "11011100";
            when "10010100" => OUTPUT <= "00100010";
            when "10010101" => OUTPUT <= "00101010";
            when "10010110" => OUTPUT <= "10010000";
            when "10010111" => OUTPUT <= "10001000";
            when "10011000" => OUTPUT <= "01000110";
            when "10011001" => OUTPUT <= "11101110";
            when "10011010" => OUTPUT <= "10111000";
            when "10011011" => OUTPUT <= "00010100";
            when "10011100" => OUTPUT <= "11011110";
            when "10011101" => OUTPUT <= "01011110";
            when "10011110" => OUTPUT <= "00001011";
            when "10011111" => OUTPUT <= "11011011";
            when "10100000" => OUTPUT <= "11100000";
            when "10100001" => OUTPUT <= "00110010";
            when "10100010" => OUTPUT <= "00111010";
            when "10100011" => OUTPUT <= "00001010";
            when "10100100" => OUTPUT <= "01001001";
            when "10100101" => OUTPUT <= "00000110";
            when "10100110" => OUTPUT <= "00100100";
            when "10100111" => OUTPUT <= "01011100";
            when "10101000" => OUTPUT <= "11000010";
            when "10101001" => OUTPUT <= "11010011";
            when "10101010" => OUTPUT <= "10101100";
            when "10101011" => OUTPUT <= "01100010";
            when "10101100" => OUTPUT <= "10010001";
            when "10101101" => OUTPUT <= "10010101";
            when "10101110" => OUTPUT <= "11100100";
            when "10101111" => OUTPUT <= "01111001";
            when "10110000" => OUTPUT <= "11100111";
            when "10110001" => OUTPUT <= "11001000";
            when "10110010" => OUTPUT <= "00110111";
            when "10110011" => OUTPUT <= "01101101";
            when "10110100" => OUTPUT <= "10001101";
            when "10110101" => OUTPUT <= "11010101";
            when "10110110" => OUTPUT <= "01001110";
            when "10110111" => OUTPUT <= "10101001";
            when "10111000" => OUTPUT <= "01101100";
            when "10111001" => OUTPUT <= "01010110";
            when "10111010" => OUTPUT <= "11110100";
            when "10111011" => OUTPUT <= "11101010";
            when "10111100" => OUTPUT <= "01100101";
            when "10111101" => OUTPUT <= "01111010";
            when "10111110" => OUTPUT <= "10101110";
            when "10111111" => OUTPUT <= "00001000";
            when "11000000" => OUTPUT <= "10111010";
            when "11000001" => OUTPUT <= "01111000";
            when "11000010" => OUTPUT <= "00100101";
            when "11000011" => OUTPUT <= "00101110";
            when "11000100" => OUTPUT <= "00011100";
            when "11000101" => OUTPUT <= "10100110";
            when "11000110" => OUTPUT <= "10110100";
            when "11000111" => OUTPUT <= "11000110";
            when "11001000" => OUTPUT <= "11101000";
            when "11001001" => OUTPUT <= "11011101";
            when "11001010" => OUTPUT <= "01110100";
            when "11001011" => OUTPUT <= "00011111";
            when "11001100" => OUTPUT <= "01001011";
            when "11001101" => OUTPUT <= "10111101";
            when "11001110" => OUTPUT <= "10001011";
            when "11001111" => OUTPUT <= "10001010";
            when "11010000" => OUTPUT <= "01110000";
            when "11010001" => OUTPUT <= "00111110";
            when "11010010" => OUTPUT <= "10110101";
            when "11010011" => OUTPUT <= "01100110";
            when "11010100" => OUTPUT <= "01001000";
            when "11010101" => OUTPUT <= "00000011";
            when "11010110" => OUTPUT <= "11110110";
            when "11010111" => OUTPUT <= "00001110";
            when "11011000" => OUTPUT <= "01100001";
            when "11011001" => OUTPUT <= "00110101";
            when "11011010" => OUTPUT <= "01010111";
            when "11011011" => OUTPUT <= "10111001";
            when "11011100" => OUTPUT <= "10000110";
            when "11011101" => OUTPUT <= "11000001";
            when "11011110" => OUTPUT <= "00011101";
            when "11011111" => OUTPUT <= "10011110";
            when "11100000" => OUTPUT <= "11100001";
            when "11100001" => OUTPUT <= "11111000";
            when "11100010" => OUTPUT <= "10011000";
            when "11100011" => OUTPUT <= "00010001";
            when "11100100" => OUTPUT <= "01101001";
            when "11100101" => OUTPUT <= "11011001";
            when "11100110" => OUTPUT <= "10001110";
            when "11100111" => OUTPUT <= "10010100";
            when "11101000" => OUTPUT <= "10011011";
            when "11101001" => OUTPUT <= "00011110";
            when "11101010" => OUTPUT <= "10000111";
            when "11101011" => OUTPUT <= "11101001";
            when "11101100" => OUTPUT <= "11001110";
            when "11101101" => OUTPUT <= "01010101";
            when "11101110" => OUTPUT <= "00101000";
            when "11101111" => OUTPUT <= "11011111";
            when "11110000" => OUTPUT <= "10001100";
            when "11110001" => OUTPUT <= "10100001";
            when "11110010" => OUTPUT <= "10001001";
            when "11110011" => OUTPUT <= "00001101";
            when "11110100" => OUTPUT <= "10111111";
            when "11110101" => OUTPUT <= "11100110";
            when "11110110" => OUTPUT <= "01000010";
            when "11110111" => OUTPUT <= "01101000";
            when "11111000" => OUTPUT <= "01000001";
            when "11111001" => OUTPUT <= "10011001";
            when "11111010" => OUTPUT <= "00101101";
            when "11111011" => OUTPUT <= "00001111";
            when "11111100" => OUTPUT <= "10110000";
            when "11111101" => OUTPUT <= "01010100";
            when "11111110" => OUTPUT <= "10111011";
            when "11111111" => OUTPUT <= "00010110";
            when others => OUTPUT <= "00000000"; -- this will never be called
        end case;
    end process;
end SBox_architecture;
